module multiplicador(a,b,c,d,e,f,g,h , o0,o1,o2,o3,o4,o5,o6,o7);

    input a,b,c,d,e,f,g,h;
    output o0,o1,o2,o3,o4,o5,o6,o7;
    wire Na,Nb,Nc,Nd,Ne,Nf,Ng,Nh;

    not not_a(Na,a);
    not not_b(Nb,b);
    not not_c(Nc,c);
    not not_d(Nd,d);
    not not_e(Ne,e);
    not not_f(Nf,f);
    not not_g(Ng,g);
    not not_h(Nh,h);

    wire o00,o01,o02,o03,o04,o05,o06,o07,o08;
    and and_o00 (o00,a,b,c,Nd,e,Nf,g);
    and and_o01 (o01,a,b,e,Nf,g,h);
    and and_o02 (o02,a,b,c,d,e,h);
    and and_o03 (o03,a,d,e,f,g,h);
    and and_o04 (o04,a,c,d,e,f);
    and and_o05 (o05,a,b,d,e,g);
    and and_o06 (o06,a,c,e,f,h);
    and and_o07 (o07,a,c,e,f,g);
    and and_o08 (o08,a,b,e,f);
    or or_o0 (o0,o00,o01,o02,o03,o04,o05,o06,o07,o08);

    wire o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,o110,o111,o112,o113,o114,o115,o116,o117,o118,o119,o120,o121,o122;
    and and_o10 (o10,a,Nb,c,Nd,e,f,Ng,Nh);
    and and_o11 (o11,a,Nc,Nd,e,Nf,g,Nh);
    and and_o12 (o12,a,Nc,d,e,Nf,Ng,h);
    and and_o13 (o13,a,b,Nc,Ne,f,g,Nh);
    and and_o14 (o14,a,b,Nc,Ne,f,g,h);
    and and_o15 (o15,a,b,Nd,e,Nf,Ng,h);
    and and_o16 (o16,a,Nb,Nc,e,f,Ng);
    and and_o17 (o17,a,b,e,Nf,Ng,Nh);
    and and_o18 (o18,a,Nb,Nc,Nd,e,g);
    and and_o19 (o19,a,Nb,Nc,e,g,Nh);
    and and_o110 (o110,a,b,d,Ne,f,h);
    and and_o111 (o111,Na,b,d,e,f,h);
    and and_o112 (o112,Na,b,c,d,e,g);
    and and_o113 (o113,a,c,d,Ne,f,g);
    and and_o114 (o114,Na,b,d,e,f,g);
    and and_o115 (o115,a,b,c,Ne,f,h);
    and and_o116 (o116,Na,b,c,e,g,h);
    and and_o117 (o117,a,c,Ne,f,g,h);
    and and_o118 (o118,a,b,c,d,f,h);
    and and_o119 (o119,a,b,d,f,g,h);
    and and_o120 (o120,Na,b,c,e,f);
    and and_o121 (o121,a,b,c,f,g);
    and and_o122 (o122,a,Nb,e,Nf);
    or or_o1 (o1,o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,o110,o111,o112,o113,o114,o115,o116,o117,o118,o119,o120,o121,o122);

    wire o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,o210,o211,o212,o213,o214,o215,o216,o217,o218,o219,o220,o221,o222,o223,o224,o225,o226,o227,o228,o229,o230,o231,o232,o233,o234;
    and and_o20 (o20,a,Nb,c,Nd,e,f,Ng,Nh);
    and and_o21 (o21,Na,b,c,Nd,e,Nf,g,Nh);
    and and_o22 (o22,a,Nc,Nd,Ne,f,Ng,h);
    and and_o23 (o23,a,Nb,Nd,Ne,f,g,Nh);
    and and_o24 (o24,a,Nb,c,d,e,Nf,h);
    and and_o25 (o25,a,b,Nc,d,e,Ng,h);
    and and_o26 (o26,a,Nb,d,e,Nf,g,h);
    and and_o27 (o27,Na,b,c,d,Ne,f,h);
    and and_o28 (o28,a,Nc,e,f,g,Nh);
    and and_o29 (o29,Na,b,d,Ne,f,g,h);
    and and_o210 (o210,Na,b,Nc,d,e,Nf,g);
    and and_o211 (o211,a,Nb,c,Ne,f,Ng,h);
    and and_o212 (o212,Na,b,Nc,e,Ng,Nh);
    and and_o213 (o213,a,b,Nd,e,Nf,Ng,h);
    and and_o214 (o214,b,Nc,Nd,e,f,g,h);
    and and_o215 (o215,Na,Nb,c,d,e,f);
    and and_o216 (o216,a,Nb,Nc,e,f,Ng);
    and and_o217 (o217,a,b,c,Nd,e,Ng);
    and and_o218 (o218,a,b,e,Nf,Ng,Nh);
    and and_o219 (o219,a,b,c,f,Ng,Nh);
    and and_o220 (o220,a,Nb,c,e,Nf,g);
    and and_o221 (o221,a,b,Ne,Nf,g,h);
    and and_o222 (o222,Na,b,c,Ne,f,g);
    and and_o223 (o223,a,Nb,Nc,Nd,f,h);
    and and_o224 (o224,b,Nc,Nd,e,g,Nh);
    and and_o225 (o225,a,Nb,Nc,Ne,f,h);
    and and_o226 (o226,a,Nb,Nc,f,g,Nh);
    and and_o227 (o227,Nb,c,d,e,g,h);
    and and_o228 (o228,a,c,d,Nf,g,h);
    and and_o229 (o229,Na,c,d,e,f,g);
    and and_o230 (o230,b,c,Ne,f,g,h);
    and and_o231 (o231,Na,b,Nc,Nd,e);
    and and_o232 (o232,Na,b,e,Nf,Ng);
    and and_o233 (o233,c,d,e,f,g,h);
    and and_o234 (o234,a,Ne,f,Ng,Nh);
    or or_o2 (o2,o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,o210,o211,o212,o213,o214,o215,o216,o217,o218,o219,o220,o221,o222,o223,o224,o225,o226,o227,o228,o229,o230,o231,o232,o233,o234);

    wire o30,o31,o32,o33,o34,o35,o36,o37,o38,o39,o310,o311,o312,o313,o314,o315,o316,o317,o318,o319,o320,o321,o322,o323,o324,o325,o326,o327,o328,o329,o330,o331,o332,o333,o334,o335,o336,o337,o338;
    and and_o30 (o30,Na,b,Nc,d,Ne,f,Ng,h);
    and and_o31 (o31,a,Nb,c,Nd,e,f,Ng,Nh);
    and and_o32 (o32,a,Nb,Nd,Ne,Nf,g);
    and and_o33 (o33,Na,b,c,Nd,e,Nf,g,Nh);
    and and_o34 (o34,a,Nb,c,d,e,Nf,g,h);
    and and_o35 (o35,a,Nb,Nc,d,e,Ng,h);
    and and_o36 (o36,Na,Nb,c,d,Ne,f,g);
    and and_o37 (o37,a,Nc,Nd,e,Nf,g,Nh);
    and and_o38 (o38,Na,b,c,Ne,Nf,g,h);
    and and_o39 (o39,a,Nb,Nd,Ne,f,g,Nh);
    and and_o310 (o310,a,Nc,d,e,Nf,Ng,h);
    and and_o311 (o311,Na,b,c,d,e,Ng);
    and and_o312 (o312,Na,c,d,Ne,f,g,h);
    and and_o313 (o313,Na,b,Nc,d,e,Nf,g);
    and and_o314 (o314,a,Nb,c,Ne,f,Ng,h);
    and and_o315 (o315,Na,Nb,c,e,Nf,Nh);
    and and_o316 (o316,Na,b,Nd,Ne,f,Ng);
    and and_o317 (o317,Na,b,Nc,Ne,f,Nh);
    and and_o318 (o318,a,b,Nc,Ne,f,g,h);
    and and_o319 (o319,b,Nc,Nd,e,f,g,h);
    and and_o320 (o320,Na,c,e,Nf,Ng);
    and and_o321 (o321,Na,b,Nc,Nd,f);
    and and_o322 (o322,a,Nb,Nc,Nd,e,g);
    and and_o323 (o323,a,Nb,Nc,e,g,Nh);
    and and_o324 (o324,a,b,c,Ne,g,Nh);
    and and_o325 (o325,Na,c,Nd,e,f,g);
    and and_o326 (o326,c,d,e,Nf,Ng,Nh);
    and and_o327 (o327,a,Nb,Nc,f,g,Nh);
    and and_o328 (o328,a,Nb,Nc,Ne,g,h);
    and and_o329 (o329,a,b,c,d,g,Nh);
    and and_o330 (o330,a,b,c,Nd,e,h);
    and and_o331 (o331,a,d,e,f,g,Nh);
    and and_o332 (o332,c,Nd,e,f,g,h);
    and and_o333 (o333,b,Nc,Nd,f,Ng);
    and and_o334 (o334,c,Nd,e,Nf,Ng);
    and and_o335 (o335,Na,Nb,c,Nd,e);
    and and_o336 (o336,b,Ne,f,Ng,Nh);
    and and_o337 (o337,a,Ne,Nf,g,Nh);
    and and_o338 (o338,b,d,f,Ng,Nh);
    or or_o3 (o3,o30,o31,o32,o33,o34,o35,o36,o37,o38,o39,o310,o311,o312,o313,o314,o315,o316,o317,o318,o319,o320,o321,o322,o323,o324,o325,o326,o327,o328,o329,o330,o331,o332,o333,o334,o335,o336,o337,o338);

    wire o40,o41,o42,o43,o44,o45,o46,o47,o48,o49,o410,o411,o412,o413,o414,o415,o416,o417,o418,o419,o420,o421,o422,o423,o424,o425,o426,o427,o428,o429,o430,o431,o432,o433,o434,o435;
    and and_o40 (o40,Na,Nb,c,d,Ne,Nf,g,h);
    and and_o41 (o41,Na,b,Nc,d,Ne,f,Ng,h);
    and and_o42 (o42,a,Nb,c,d,e,f,Ng,h);
    and and_o43 (o43,a,b,Nc,d,e,Nf,g,h);
    and and_o44 (o44,Na,b,c,Nd,e,Nf,g,Nh);
    and and_o45 (o45,a,Nb,c,d,e,Nf,g,h);
    and and_o46 (o46,a,Nc,Nd,Ne,f,Ng,h);
    and and_o47 (o47,a,b,Nc,e,f,Ng,h);
    and and_o48 (o48,a,b,Nc,Ne,f,g,Nh);
    and and_o49 (o49,a,b,c,Nd,e,Nf,g);
    and and_o410 (o410,Na,Nb,c,Ne,f,Ng);
    and and_o411 (o411,Na,b,Nc,Ne,Nf,g);
    and and_o412 (o412,a,b,Nd,e,Nf,Ng,h);
    and and_o413 (o413,a,b,c,Ne,Nf,h);
    and and_o414 (o414,a,Nb,Nc,Nd,f,h);
    and and_o415 (o415,c,d,e,Nf,Ng,Nh);
    and and_o416 (o416,b,Nc,Nd,e,g,Nh);
    and and_o417 (o417,a,Nb,Nc,Ne,f,h);
    and and_o418 (o418,a,Nb,Nc,Ne,g,h);
    and and_o419 (o419,a,b,c,d,Ne,h);
    and and_o420 (o420,Na,b,c,d,e,h);
    and and_o421 (o421,a,d,Ne,f,g,h);
    and and_o422 (o422,Na,d,e,f,g,h);
    and and_o423 (o423,a,Nb,Nd,Nf,h);
    and and_o424 (o424,Nb,c,Nd,f,Nh);
    and and_o425 (o425,Na,Nb,Nc,d,e);
    and and_o426 (o426,Nc,d,e,Ng,Nh);
    and and_o427 (o427,c,Nd,f,Ng,Nh);
    and and_o428 (o428,Na,d,e,Nf,Ng);
    and and_o429 (o429,Na,b,Nc,Nd,g);
    and and_o430 (o430,a,Ne,Nf,Ng,h);
    and and_o431 (o431,c,Ne,f,Ng,Nh);
    and and_o432 (o432,b,Ne,Nf,g,Nh);
    and and_o433 (o433,Nb,d,e,g,Nh);
    and and_o434 (o434,b,d,Ne,g,Nh);
    and and_o435 (o435,Na,c,Nd,f,h);
    or or_o4 (o4,o40,o41,o42,o43,o44,o45,o46,o47,o48,o49,o410,o411,o412,o413,o414,o415,o416,o417,o418,o419,o420,o421,o422,o423,o424,o425,o426,o427,o428,o429,o430,o431,o432,o433,o434,o435);

    wire o50,o51,o52,o53,o54,o55,o56,o57,o58;
    and and_o50 (o50,Nc,d,f,Nh);
    and and_o51 (o51,b,Nc,Nd,h);
    and and_o52 (o52,d,f,Ng,Nh);
    and and_o53 (o53,b,Nd,Ng,h);
    and and_o54 (o54,Nb,c,Nd,g);
    and and_o55 (o55,c,Nd,g,Nh);
    and and_o56 (o56,c,Nf,g,Nh);
    and and_o57 (o57,b,d,Nf,h);
    and and_o58 (o58,Nb,d,f,h);
    or or_o5 (o5,o50,o51,o52,o53,o54,o55,o56,o57,o58);

    wire o60,o61,o62,o63;
    and and_o60 (o60,c,Nd,h);
    and and_o61 (o61,Nc,d,g);
    and and_o62 (o62,d,g,Nh);
    and and_o63 (o63,c,Ng,h);
    or or_o6 (o6,o60,o61,o62,o63);

    wire o70;
    and and_o70 (o70,d,h);
    or or_o7 (o7,o70);

endmodule
